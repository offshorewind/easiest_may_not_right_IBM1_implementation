ställ konen på den röda kvadraten på kvadraten
ta konen på kvadraten
ta blocket
ställ den röda konen på kvadraten
ställ blocket på den blåa kvadraten på kvadraten
ställ den gröna konen på den blåa cirkeln
ställ den gröna konen på den röda kvadraten
ställ det blåa blocket på den röda kvadraten
ställ det röda blocket på den röda kvadraten
ställ den röda konen på den gröna cirkeln på kvadraten
ta den gröna kuben på den röda cirkeln
ta den blåa kuben på den gröna cirkeln
ställ blocket på cirkeln på den röda kvadraten
ta kuben
ta blocket
ställ blocket på cirkeln på kvadraten
ta det gröna blocket
ta kuben på den röda cirkeln
ställ blocket på den röda kvadraten
ställ blocket på kvadraten på den röda cirkeln
ta kuben
ställ den röda konen på kvadraten
ställ kuben på cirkeln på den röda cirkeln
ställ det blåa blocket på den blåa kvadraten
ta blocket på kvadraten
ta det röda blocket
ta den röda kuben på kvadraten
ställ konen på den röda kvadraten på den röda kvadraten
ställ blocket på den röda cirkeln
ta det gröna blocket
ställ blocket på den röda cirkeln
ställ den blåa kuben på den röda kvadraten
ställ det blåa blocket på den blåa kvadraten
ta konen
ställ konen på den röda cirkeln på kvadraten
ta det gröna blocket
ställ konen på kvadraten på den röda kvadraten
ställ kuben på kvadraten på cirkeln
ta blocket på den röda cirkeln
ta blocket
ställ den röda kuben på den röda kvadraten
ta det blåa blocket
ta blocket
ta det gröna blocket
ställ den blåa kuben på kvadraten
ställ blocket på kvadraten på den blåa cirkeln
ställ kuben på den röda cirkeln på den röda kvadraten
ta det röda blocket
ställ den blåa kuben på den gröna cirkeln
ställ det röda blocket på den blåa cirkeln
ställ kuben på kvadraten
ställ den blåa konen på kvadraten på kvadraten
ställ konen på den röda cirkeln på kvadraten
ställ det blåa blocket på den röda cirkeln
ställ kuben på den röda cirkeln på cirkeln
ta kuben
ställ den blåa konen på cirkeln
ta konen
ställ den blåa konen på den röda cirkeln på kvadraten
ställ den röda kuben på den röda kvadraten
ställ blocket på den blåa cirkeln
ta kuben på cirkeln
ställ kuben på cirkeln på cirkeln
ställ blocket på den röda kvadraten
ta blocket på cirkeln
ställ det gröna blocket på den gröna kvadraten
ta det röda blocket
ta konen
ställ kuben på kvadraten
ta den röda konen
ställ konen på kvadraten på den röda cirkeln
ställ den röda konen på cirkeln
ställ konen på cirkeln på den röda cirkeln
ta det röda blocket på den blåa kvadraten
ta det röda blocket
ta blocket
ställ det röda blocket på den gröna cirkeln
ställ blocket på cirkeln på cirkeln
ställ konen på cirkeln på den röda cirkeln
ställ det röda blocket på cirkeln
ställ konen på kvadraten
ställ blocket på den blåa kvadraten på kvadraten
ställ kuben på den röda cirkeln
ta det röda blocket
ställ det röda blocket på cirkeln på den blåa kvadraten
ställ kuben på den röda kvadraten på cirkeln
ställ den blåa konen på den blåa cirkeln
ställ blocket på kvadraten
ställ kuben på cirkeln
ta det gröna blocket
ställ den röda konen på kvadraten på cirkeln
ställ blocket på den röda cirkeln
ställ den blåa konen på den röda kvadraten
ställ den röda konen på cirkeln
ställ den blåa konen på den röda cirkeln på cirkeln
ta den blåa konen
ställ det röda blocket på den gröna cirkeln
ställ det gröna blocket på den röda kvadraten
ställ kuben på den gröna kvadraten
ta det blåa blocket
